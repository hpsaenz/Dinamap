[FSV][0][Vital signs (ProCare)][Enterprise, Medicalogic][2.000000][55.000000, 61.000000, 2641.000000, 60.000000, 56.000000, 4747.000000, 57.000000, 54.000000, 53.000000, 2173.000000]
[EFS][3][Vital signs (ProCare)][Enterprise, MedicaLogic][Version 5.5_1.0 DINAMAP ProCare basic vital signs with in-line text translation; Authored at: GE Medical Systems on 9/12/2003 11:07:25 AM with 2.5.1_7][Vital Signs][VITALS.EFM][VITALS.XLT][VITALS.XLW][VITALS.PEF][][1][Arial]
