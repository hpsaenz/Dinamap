[EFS][3][Vital signs (ProCare)][Enterprise, MedicaLogic][Version 5.5_1.0 DINAMAP ProCare basic vital signs with in-line text translation; Authored at: Memorial Family Practice, Site # 196 on 10/19/2015 4:45:13 PM with 6.25][Vital Signs][VITALS.EFM][VITALS.XLT][VITALS.XLW][VITALS.PEF][][1][Arial][]